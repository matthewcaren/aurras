`timescale 1ns / 1ps
`default_nettype none

module frequency_sweep (
  input wire clk_in,
  input wire rst_in,
  output wire [15:0] sound_out
);

// Paramaters to be adjusted based on desired outcome



 

endmodule


`timescale 1ns / 1ps
`default_nettype wire
